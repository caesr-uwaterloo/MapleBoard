module test_run_elf;
  initial begin
    $display("Hello World from test_run_elf");
  end
endmodule
